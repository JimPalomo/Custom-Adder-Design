-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"
-- CREATED		"Tue Nov 10 14:33:56 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY IL_level5_new IS 
	PORT
	(
		NZFlag :  IN  STD_LOGIC;
		Cout_0 :  IN  STD_LOGIC;
		In_3 :  IN  STD_LOGIC;
		In_2 :  IN  STD_LOGIC;
		In_1 :  IN  STD_LOGIC;
		In_0 :  IN  STD_LOGIC;
		LSZD_Pos0 :  IN  STD_LOGIC;
		LSZD_Pos1 :  IN  STD_LOGIC;
		LSZD_Pos2 :  IN  STD_LOGIC;
		In_4 :  IN  STD_LOGIC;
		In_5 :  IN  STD_LOGIC;
		In_6 :  IN  STD_LOGIC;
		In_7 :  IN  STD_LOGIC;
		LSZD_Pos3 :  IN  STD_LOGIC;
		In_8 :  IN  STD_LOGIC;
		In_9 :  IN  STD_LOGIC;
		In_10 :  IN  STD_LOGIC;
		In_11 :  IN  STD_LOGIC;
		In_12 :  IN  STD_LOGIC;
		In_13 :  IN  STD_LOGIC;
		In_14 :  IN  STD_LOGIC;
		In_15 :  IN  STD_LOGIC;
		LSZD_Pos4 :  IN  STD_LOGIC;
		In_16 :  IN  STD_LOGIC;
		In_17 :  IN  STD_LOGIC;
		In_18 :  IN  STD_LOGIC;
		In_19 :  IN  STD_LOGIC;
		In_20 :  IN  STD_LOGIC;
		In_21 :  IN  STD_LOGIC;
		In_22 :  IN  STD_LOGIC;
		In_23 :  IN  STD_LOGIC;
		In_24 :  IN  STD_LOGIC;
		In_25 :  IN  STD_LOGIC;
		In_26 :  IN  STD_LOGIC;
		In_27 :  IN  STD_LOGIC;
		In_28 :  IN  STD_LOGIC;
		In_29 :  IN  STD_LOGIC;
		In_30 :  IN  STD_LOGIC;
		In_31 :  IN  STD_LOGIC;
		LSZD_Pos5 :  IN  STD_LOGIC;
		In_32 :  IN  STD_LOGIC;
		Out_3 :  OUT  STD_LOGIC;
		Out_2 :  OUT  STD_LOGIC;
		Out_1 :  OUT  STD_LOGIC;
		Out_0 :  OUT  STD_LOGIC;
		Out_4 :  OUT  STD_LOGIC;
		Out_5 :  OUT  STD_LOGIC;
		Out_6 :  OUT  STD_LOGIC;
		Out_7 :  OUT  STD_LOGIC;
		Out_28 :  OUT  STD_LOGIC;
		Out_8 :  OUT  STD_LOGIC;
		Out_9 :  OUT  STD_LOGIC;
		Out_11 :  OUT  STD_LOGIC;
		Out_10 :  OUT  STD_LOGIC;
		Out_12 :  OUT  STD_LOGIC;
		Out_13 :  OUT  STD_LOGIC;
		Out_14 :  OUT  STD_LOGIC;
		Out_15 :  OUT  STD_LOGIC;
		Out_16 :  OUT  STD_LOGIC;
		Out_17 :  OUT  STD_LOGIC;
		Out_18 :  OUT  STD_LOGIC;
		Out_19 :  OUT  STD_LOGIC;
		Out_20 :  OUT  STD_LOGIC;
		Out_21 :  OUT  STD_LOGIC;
		Out_22 :  OUT  STD_LOGIC;
		Out_23 :  OUT  STD_LOGIC;
		Out_24 :  OUT  STD_LOGIC;
		Out_25 :  OUT  STD_LOGIC;
		Out_26 :  OUT  STD_LOGIC;
		Out_27 :  OUT  STD_LOGIC;
		Out_29 :  OUT  STD_LOGIC;
		Out_30 :  OUT  STD_LOGIC;
		Out_31 :  OUT  STD_LOGIC;
		Out_32 :  OUT  STD_LOGIC
	);
END IL_level5_new;

ARCHITECTURE bdf_type OF IL_level5_new IS 

COMPONENT decoder6_64
	PORT(i0 : IN STD_LOGIC;
		 i1 : IN STD_LOGIC;
		 i2 : IN STD_LOGIC;
		 i3 : IN STD_LOGIC;
		 i4 : IN STD_LOGIC;
		 i5 : IN STD_LOGIC;
		 En : IN STD_LOGIC;
		 d0 : OUT STD_LOGIC;
		 d1 : OUT STD_LOGIC;
		 d2 : OUT STD_LOGIC;
		 d3 : OUT STD_LOGIC;
		 d4 : OUT STD_LOGIC;
		 d5 : OUT STD_LOGIC;
		 d6 : OUT STD_LOGIC;
		 d7 : OUT STD_LOGIC;
		 d8 : OUT STD_LOGIC;
		 d9 : OUT STD_LOGIC;
		 d10 : OUT STD_LOGIC;
		 d11 : OUT STD_LOGIC;
		 d12 : OUT STD_LOGIC;
		 d13 : OUT STD_LOGIC;
		 d14 : OUT STD_LOGIC;
		 d15 : OUT STD_LOGIC;
		 d16 : OUT STD_LOGIC;
		 d17 : OUT STD_LOGIC;
		 d18 : OUT STD_LOGIC;
		 d19 : OUT STD_LOGIC;
		 d20 : OUT STD_LOGIC;
		 d21 : OUT STD_LOGIC;
		 d22 : OUT STD_LOGIC;
		 d23 : OUT STD_LOGIC;
		 d24 : OUT STD_LOGIC;
		 d25 : OUT STD_LOGIC;
		 d26 : OUT STD_LOGIC;
		 d27 : OUT STD_LOGIC;
		 d28 : OUT STD_LOGIC;
		 d29 : OUT STD_LOGIC;
		 d30 : OUT STD_LOGIC;
		 d31 : OUT STD_LOGIC;
		 d32 : OUT STD_LOGIC;
		 d33 : OUT STD_LOGIC;
		 d34 : OUT STD_LOGIC;
		 d35 : OUT STD_LOGIC;
		 d36 : OUT STD_LOGIC;
		 d37 : OUT STD_LOGIC;
		 d38 : OUT STD_LOGIC;
		 d39 : OUT STD_LOGIC;
		 d40 : OUT STD_LOGIC;
		 d41 : OUT STD_LOGIC;
		 d42 : OUT STD_LOGIC;
		 d43 : OUT STD_LOGIC;
		 d44 : OUT STD_LOGIC;
		 d45 : OUT STD_LOGIC;
		 d46 : OUT STD_LOGIC;
		 d47 : OUT STD_LOGIC;
		 d48 : OUT STD_LOGIC;
		 d49 : OUT STD_LOGIC;
		 d50 : OUT STD_LOGIC;
		 d51 : OUT STD_LOGIC;
		 d52 : OUT STD_LOGIC;
		 d53 : OUT STD_LOGIC;
		 d54 : OUT STD_LOGIC;
		 d55 : OUT STD_LOGIC;
		 d56 : OUT STD_LOGIC;
		 d57 : OUT STD_LOGIC;
		 d58 : OUT STD_LOGIC;
		 d59 : OUT STD_LOGIC;
		 d60 : OUT STD_LOGIC;
		 d61 : OUT STD_LOGIC;
		 d62 : OUT STD_LOGIC;
		 d63 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mux2_1
	PORT(I_0 : IN STD_LOGIC;
		 Sel : IN STD_LOGIC;
		 I_1 : IN STD_LOGIC;
		 Out_0 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;


BEGIN 



b2v_inst1 : decoder6_64
PORT MAP(i0 => LSZD_Pos0,
		 i1 => LSZD_Pos1,
		 i2 => LSZD_Pos2,
		 i3 => LSZD_Pos3,
		 i4 => LSZD_Pos4,
		 i5 => LSZD_Pos5,
		 En => SYNTHESIZED_WIRE_0,
		 d0 => SYNTHESIZED_WIRE_68,
		 d1 => SYNTHESIZED_WIRE_54,
		 d2 => SYNTHESIZED_WIRE_22,
		 d3 => SYNTHESIZED_WIRE_4,
		 d4 => SYNTHESIZED_WIRE_6,
		 d5 => SYNTHESIZED_WIRE_18,
		 d6 => SYNTHESIZED_WIRE_20,
		 d7 => SYNTHESIZED_WIRE_32,
		 d8 => SYNTHESIZED_WIRE_34,
		 d9 => SYNTHESIZED_WIRE_36,
		 d10 => SYNTHESIZED_WIRE_40,
		 d11 => SYNTHESIZED_WIRE_42,
		 d12 => SYNTHESIZED_WIRE_44,
		 d13 => SYNTHESIZED_WIRE_46,
		 d14 => SYNTHESIZED_WIRE_48,
		 d15 => SYNTHESIZED_WIRE_70,
		 d16 => SYNTHESIZED_WIRE_66,
		 d17 => SYNTHESIZED_WIRE_38,
		 d18 => SYNTHESIZED_WIRE_74,
		 d19 => SYNTHESIZED_WIRE_76,
		 d20 => SYNTHESIZED_WIRE_78,
		 d21 => SYNTHESIZED_WIRE_80,
		 d22 => SYNTHESIZED_WIRE_82,
		 d23 => SYNTHESIZED_WIRE_84,
		 d24 => SYNTHESIZED_WIRE_86,
		 d25 => SYNTHESIZED_WIRE_88,
		 d26 => SYNTHESIZED_WIRE_90,
		 d27 => SYNTHESIZED_WIRE_92,
		 d28 => SYNTHESIZED_WIRE_94,
		 d29 => SYNTHESIZED_WIRE_96,
		 d30 => SYNTHESIZED_WIRE_131,
		 d31 => SYNTHESIZED_WIRE_10,
		 d32 => SYNTHESIZED_WIRE_132);


SYNTHESIZED_WIRE_121 <= NOT(NZFlag);



SYNTHESIZED_WIRE_2 <= NOT(In_32);



b2v_inst103 : mux2_1
PORT MAP(I_0 => In_32,
		 Sel => SYNTHESIZED_WIRE_132,
		 I_1 => SYNTHESIZED_WIRE_2,
		 Out_0 => Out_32);


SYNTHESIZED_WIRE_14 <= NOT(In_1);



SYNTHESIZED_WIRE_16 <= NOT(In_0);



SYNTHESIZED_WIRE_135 <= SYNTHESIZED_WIRE_133 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_133 <= SYNTHESIZED_WIRE_134 OR SYNTHESIZED_WIRE_6;


b2v_inst162 : mux2_1
PORT MAP(I_0 => In_3,
		 Sel => SYNTHESIZED_WIRE_135,
		 I_1 => SYNTHESIZED_WIRE_8,
		 Out_0 => Out_3);


SYNTHESIZED_WIRE_163 <= SYNTHESIZED_WIRE_132 OR SYNTHESIZED_WIRE_10;


b2v_inst165 : mux2_1
PORT MAP(I_0 => In_2,
		 Sel => SYNTHESIZED_WIRE_136,
		 I_1 => SYNTHESIZED_WIRE_12,
		 Out_0 => Out_2);


b2v_inst166 : mux2_1
PORT MAP(I_0 => In_1,
		 Sel => SYNTHESIZED_WIRE_137,
		 I_1 => SYNTHESIZED_WIRE_14,
		 Out_0 => Out_1);


b2v_inst167 : mux2_1
PORT MAP(I_0 => In_0,
		 Sel => SYNTHESIZED_WIRE_15,
		 I_1 => SYNTHESIZED_WIRE_16,
		 Out_0 => Out_0);


SYNTHESIZED_WIRE_134 <= SYNTHESIZED_WIRE_138 OR SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_138 <= SYNTHESIZED_WIRE_139 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_24 <= NOT(In_4);



SYNTHESIZED_WIRE_136 <= SYNTHESIZED_WIRE_135 OR SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_26 <= NOT(In_5);



b2v_inst21 : mux2_1
PORT MAP(I_0 => In_4,
		 Sel => SYNTHESIZED_WIRE_133,
		 I_1 => SYNTHESIZED_WIRE_24,
		 Out_0 => Out_4);


b2v_inst22 : mux2_1
PORT MAP(I_0 => In_5,
		 Sel => SYNTHESIZED_WIRE_134,
		 I_1 => SYNTHESIZED_WIRE_26,
		 Out_0 => Out_5);


SYNTHESIZED_WIRE_28 <= NOT(In_6);



b2v_inst24 : mux2_1
PORT MAP(I_0 => In_6,
		 Sel => SYNTHESIZED_WIRE_138,
		 I_1 => SYNTHESIZED_WIRE_28,
		 Out_0 => Out_6);


SYNTHESIZED_WIRE_30 <= NOT(In_7);



b2v_inst26 : mux2_1
PORT MAP(I_0 => In_7,
		 Sel => SYNTHESIZED_WIRE_139,
		 I_1 => SYNTHESIZED_WIRE_30,
		 Out_0 => Out_7);


SYNTHESIZED_WIRE_139 <= SYNTHESIZED_WIRE_140 OR SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_140 <= SYNTHESIZED_WIRE_141 OR SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_141 <= SYNTHESIZED_WIRE_142 OR SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_149 <= SYNTHESIZED_WIRE_143 OR SYNTHESIZED_WIRE_38;


SYNTHESIZED_WIRE_142 <= SYNTHESIZED_WIRE_144 OR SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_144 <= SYNTHESIZED_WIRE_145 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_145 <= SYNTHESIZED_WIRE_146 OR SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_146 <= SYNTHESIZED_WIRE_147 OR SYNTHESIZED_WIRE_46;


SYNTHESIZED_WIRE_147 <= SYNTHESIZED_WIRE_148 OR SYNTHESIZED_WIRE_48;


SYNTHESIZED_WIRE_50 <= NOT(In_9);



b2v_inst36 : mux2_1
PORT MAP(I_0 => In_9,
		 Sel => SYNTHESIZED_WIRE_141,
		 I_1 => SYNTHESIZED_WIRE_50,
		 Out_0 => Out_9);


SYNTHESIZED_WIRE_52 <= NOT(In_10);



b2v_inst38 : mux2_1
PORT MAP(I_0 => In_10,
		 Sel => SYNTHESIZED_WIRE_142,
		 I_1 => SYNTHESIZED_WIRE_52,
		 Out_0 => Out_10);


SYNTHESIZED_WIRE_56 <= NOT(In_8);



SYNTHESIZED_WIRE_137 <= SYNTHESIZED_WIRE_136 OR SYNTHESIZED_WIRE_54;


b2v_inst40 : mux2_1
PORT MAP(I_0 => In_8,
		 Sel => SYNTHESIZED_WIRE_140,
		 I_1 => SYNTHESIZED_WIRE_56,
		 Out_0 => Out_8);


SYNTHESIZED_WIRE_58 <= NOT(In_12);



b2v_inst42 : mux2_1
PORT MAP(I_0 => In_12,
		 Sel => SYNTHESIZED_WIRE_145,
		 I_1 => SYNTHESIZED_WIRE_58,
		 Out_0 => Out_12);


SYNTHESIZED_WIRE_60 <= NOT(In_13);



b2v_inst44 : mux2_1
PORT MAP(I_0 => In_13,
		 Sel => SYNTHESIZED_WIRE_146,
		 I_1 => SYNTHESIZED_WIRE_60,
		 Out_0 => Out_13);


SYNTHESIZED_WIRE_62 <= NOT(In_11);



b2v_inst46 : mux2_1
PORT MAP(I_0 => In_11,
		 Sel => SYNTHESIZED_WIRE_144,
		 I_1 => SYNTHESIZED_WIRE_62,
		 Out_0 => Out_11);


SYNTHESIZED_WIRE_64 <= NOT(In_15);



b2v_inst48 : mux2_1
PORT MAP(I_0 => In_15,
		 Sel => SYNTHESIZED_WIRE_148,
		 I_1 => SYNTHESIZED_WIRE_64,
		 Out_0 => Out_15);


SYNTHESIZED_WIRE_150 <= SYNTHESIZED_WIRE_149 OR SYNTHESIZED_WIRE_66;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_137 OR SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_148 <= SYNTHESIZED_WIRE_150 OR SYNTHESIZED_WIRE_70;


SYNTHESIZED_WIRE_72 <= NOT(In_14);



b2v_inst52 : mux2_1
PORT MAP(I_0 => In_14,
		 Sel => SYNTHESIZED_WIRE_147,
		 I_1 => SYNTHESIZED_WIRE_72,
		 Out_0 => Out_14);


SYNTHESIZED_WIRE_143 <= SYNTHESIZED_WIRE_151 OR SYNTHESIZED_WIRE_74;


SYNTHESIZED_WIRE_151 <= SYNTHESIZED_WIRE_152 OR SYNTHESIZED_WIRE_76;


SYNTHESIZED_WIRE_152 <= SYNTHESIZED_WIRE_153 OR SYNTHESIZED_WIRE_78;


SYNTHESIZED_WIRE_153 <= SYNTHESIZED_WIRE_154 OR SYNTHESIZED_WIRE_80;


SYNTHESIZED_WIRE_154 <= SYNTHESIZED_WIRE_155 OR SYNTHESIZED_WIRE_82;


SYNTHESIZED_WIRE_155 <= SYNTHESIZED_WIRE_156 OR SYNTHESIZED_WIRE_84;


SYNTHESIZED_WIRE_156 <= SYNTHESIZED_WIRE_157 OR SYNTHESIZED_WIRE_86;


SYNTHESIZED_WIRE_157 <= SYNTHESIZED_WIRE_158 OR SYNTHESIZED_WIRE_88;


SYNTHESIZED_WIRE_158 <= SYNTHESIZED_WIRE_159 OR SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_159 <= SYNTHESIZED_WIRE_160 OR SYNTHESIZED_WIRE_92;


SYNTHESIZED_WIRE_160 <= SYNTHESIZED_WIRE_161 OR SYNTHESIZED_WIRE_94;


SYNTHESIZED_WIRE_161 <= SYNTHESIZED_WIRE_162 OR SYNTHESIZED_WIRE_96;


SYNTHESIZED_WIRE_98 <= NOT(In_17);



b2v_inst66 : mux2_1
PORT MAP(I_0 => In_17,
		 Sel => SYNTHESIZED_WIRE_149,
		 I_1 => SYNTHESIZED_WIRE_98,
		 Out_0 => Out_17);


SYNTHESIZED_WIRE_100 <= NOT(In_18);



b2v_inst68 : mux2_1
PORT MAP(I_0 => In_18,
		 Sel => SYNTHESIZED_WIRE_143,
		 I_1 => SYNTHESIZED_WIRE_100,
		 Out_0 => Out_18);


SYNTHESIZED_WIRE_102 <= NOT(In_16);



SYNTHESIZED_WIRE_8 <= NOT(In_3);



b2v_inst70 : mux2_1
PORT MAP(I_0 => In_16,
		 Sel => SYNTHESIZED_WIRE_150,
		 I_1 => SYNTHESIZED_WIRE_102,
		 Out_0 => Out_16);


SYNTHESIZED_WIRE_104 <= NOT(In_20);



b2v_inst72 : mux2_1
PORT MAP(I_0 => In_20,
		 Sel => SYNTHESIZED_WIRE_152,
		 I_1 => SYNTHESIZED_WIRE_104,
		 Out_0 => Out_20);


SYNTHESIZED_WIRE_106 <= NOT(In_21);



b2v_inst74 : mux2_1
PORT MAP(I_0 => In_21,
		 Sel => SYNTHESIZED_WIRE_153,
		 I_1 => SYNTHESIZED_WIRE_106,
		 Out_0 => Out_21);


SYNTHESIZED_WIRE_108 <= NOT(In_19);



b2v_inst76 : mux2_1
PORT MAP(I_0 => In_19,
		 Sel => SYNTHESIZED_WIRE_151,
		 I_1 => SYNTHESIZED_WIRE_108,
		 Out_0 => Out_19);


SYNTHESIZED_WIRE_110 <= NOT(In_23);



b2v_inst78 : mux2_1
PORT MAP(I_0 => In_23,
		 Sel => SYNTHESIZED_WIRE_155,
		 I_1 => SYNTHESIZED_WIRE_110,
		 Out_0 => Out_23);


SYNTHESIZED_WIRE_112 <= NOT(In_24);



SYNTHESIZED_WIRE_12 <= NOT(In_2);



b2v_inst80 : mux2_1
PORT MAP(I_0 => In_24,
		 Sel => SYNTHESIZED_WIRE_156,
		 I_1 => SYNTHESIZED_WIRE_112,
		 Out_0 => Out_24);


SYNTHESIZED_WIRE_114 <= NOT(In_22);



b2v_inst82 : mux2_1
PORT MAP(I_0 => In_22,
		 Sel => SYNTHESIZED_WIRE_154,
		 I_1 => SYNTHESIZED_WIRE_114,
		 Out_0 => Out_22);


SYNTHESIZED_WIRE_116 <= NOT(In_26);



b2v_inst84 : mux2_1
PORT MAP(I_0 => In_26,
		 Sel => SYNTHESIZED_WIRE_158,
		 I_1 => SYNTHESIZED_WIRE_116,
		 Out_0 => Out_26);


SYNTHESIZED_WIRE_118 <= NOT(In_27);



b2v_inst86 : mux2_1
PORT MAP(I_0 => In_27,
		 Sel => SYNTHESIZED_WIRE_159,
		 I_1 => SYNTHESIZED_WIRE_118,
		 Out_0 => Out_27);


SYNTHESIZED_WIRE_120 <= NOT(In_25);



b2v_inst88 : mux2_1
PORT MAP(I_0 => In_25,
		 Sel => SYNTHESIZED_WIRE_157,
		 I_1 => SYNTHESIZED_WIRE_120,
		 Out_0 => Out_25);


SYNTHESIZED_WIRE_123 <= NOT(In_28);



SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_121 AND Cout_0;


b2v_inst90 : mux2_1
PORT MAP(I_0 => In_28,
		 Sel => SYNTHESIZED_WIRE_160,
		 I_1 => SYNTHESIZED_WIRE_123,
		 Out_0 => Out_28);


SYNTHESIZED_WIRE_125 <= NOT(In_30);



b2v_inst92 : mux2_1
PORT MAP(I_0 => In_30,
		 Sel => SYNTHESIZED_WIRE_162,
		 I_1 => SYNTHESIZED_WIRE_125,
		 Out_0 => Out_30);


SYNTHESIZED_WIRE_127 <= NOT(In_31);



b2v_inst94 : mux2_1
PORT MAP(I_0 => In_31,
		 Sel => SYNTHESIZED_WIRE_163,
		 I_1 => SYNTHESIZED_WIRE_127,
		 Out_0 => Out_31);


SYNTHESIZED_WIRE_129 <= NOT(In_29);



b2v_inst96 : mux2_1
PORT MAP(I_0 => In_29,
		 Sel => SYNTHESIZED_WIRE_161,
		 I_1 => SYNTHESIZED_WIRE_129,
		 Out_0 => Out_29);


SYNTHESIZED_WIRE_162 <= SYNTHESIZED_WIRE_163 OR SYNTHESIZED_WIRE_131;


END bdf_type;