-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"
-- CREATED		"Tue Nov 10 15:07:29 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY ACL_adder IS 
	PORT
	(
		cin_init :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		a :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		b :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		sum :  OUT  STD_LOGIC_VECTOR(64 DOWNTO 0)
	);
END ACL_adder;

ARCHITECTURE bdf_type OF ACL_adder IS 

COMPONENT il_level5_new
	PORT(LSZD_Pos0 : IN STD_LOGIC;
		 LSZD_Pos1 : IN STD_LOGIC;
		 LSZD_Pos2 : IN STD_LOGIC;
		 LSZD_Pos3 : IN STD_LOGIC;
		 LSZD_Pos4 : IN STD_LOGIC;
		 LSZD_Pos5 : IN STD_LOGIC;
		 NZFlag : IN STD_LOGIC;
		 Cout_0 : IN STD_LOGIC;
		 In_0 : IN STD_LOGIC;
		 In_1 : IN STD_LOGIC;
		 In_2 : IN STD_LOGIC;
		 In_3 : IN STD_LOGIC;
		 In_4 : IN STD_LOGIC;
		 In_5 : IN STD_LOGIC;
		 In_6 : IN STD_LOGIC;
		 In_7 : IN STD_LOGIC;
		 In_8 : IN STD_LOGIC;
		 In_9 : IN STD_LOGIC;
		 In_10 : IN STD_LOGIC;
		 In_11 : IN STD_LOGIC;
		 In_12 : IN STD_LOGIC;
		 In_13 : IN STD_LOGIC;
		 In_14 : IN STD_LOGIC;
		 In_15 : IN STD_LOGIC;
		 In_16 : IN STD_LOGIC;
		 In_17 : IN STD_LOGIC;
		 In_18 : IN STD_LOGIC;
		 In_19 : IN STD_LOGIC;
		 In_20 : IN STD_LOGIC;
		 In_21 : IN STD_LOGIC;
		 In_22 : IN STD_LOGIC;
		 In_23 : IN STD_LOGIC;
		 In_24 : IN STD_LOGIC;
		 In_25 : IN STD_LOGIC;
		 In_26 : IN STD_LOGIC;
		 In_27 : IN STD_LOGIC;
		 In_28 : IN STD_LOGIC;
		 In_29 : IN STD_LOGIC;
		 In_30 : IN STD_LOGIC;
		 In_31 : IN STD_LOGIC;
		 In_32 : IN STD_LOGIC;
		 Out_0 : OUT STD_LOGIC;
		 Out_1 : OUT STD_LOGIC;
		 Out_2 : OUT STD_LOGIC;
		 Out_3 : OUT STD_LOGIC;
		 Out_4 : OUT STD_LOGIC;
		 Out_5 : OUT STD_LOGIC;
		 Out_6 : OUT STD_LOGIC;
		 Out_7 : OUT STD_LOGIC;
		 Out_8 : OUT STD_LOGIC;
		 Out_9 : OUT STD_LOGIC;
		 Out_10 : OUT STD_LOGIC;
		 Out_11 : OUT STD_LOGIC;
		 Out_12 : OUT STD_LOGIC;
		 Out_13 : OUT STD_LOGIC;
		 Out_14 : OUT STD_LOGIC;
		 Out_15 : OUT STD_LOGIC;
		 Out_16 : OUT STD_LOGIC;
		 Out_17 : OUT STD_LOGIC;
		 Out_18 : OUT STD_LOGIC;
		 Out_19 : OUT STD_LOGIC;
		 Out_20 : OUT STD_LOGIC;
		 Out_21 : OUT STD_LOGIC;
		 Out_22 : OUT STD_LOGIC;
		 Out_23 : OUT STD_LOGIC;
		 Out_24 : OUT STD_LOGIC;
		 Out_25 : OUT STD_LOGIC;
		 Out_26 : OUT STD_LOGIC;
		 Out_27 : OUT STD_LOGIC;
		 Out_28 : OUT STD_LOGIC;
		 Out_29 : OUT STD_LOGIC;
		 Out_30 : OUT STD_LOGIC;
		 Out_31 : OUT STD_LOGIC;
		 Out_32 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT leaf
	PORT(A_1 : IN STD_LOGIC;
		 B_1 : IN STD_LOGIC;
		 A_0 : IN STD_LOGIC;
		 B_0 : IN STD_LOGIC;
		 Sum_1p : OUT STD_LOGIC;
		 Cout_1p : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC;
		 Sum_0 : OUT STD_LOGIC;
		 Pos : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT il_level2
	PORT(LSZD_Pos0 : IN STD_LOGIC;
		 LSZD_Pos1 : IN STD_LOGIC;
		 LSZD_Pos2 : IN STD_LOGIC;
		 Cout_0 : IN STD_LOGIC;
		 In_0 : IN STD_LOGIC;
		 In_1 : IN STD_LOGIC;
		 In_2 : IN STD_LOGIC;
		 In_3 : IN STD_LOGIC;
		 In_4 : IN STD_LOGIC;
		 Out_0 : OUT STD_LOGIC;
		 Out_1 : OUT STD_LOGIC;
		 Out_2 : OUT STD_LOGIC;
		 Out_3 : OUT STD_LOGIC;
		 Out_4 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lszd_level1
	PORT(MS0 : IN STD_LOGIC;
		 MSH_LS_sumbit : IN STD_LOGIC;
		 NZ_MS : IN STD_LOGIC;
		 NZ_LS : IN STD_LOGIC;
		 P1 : OUT STD_LOGIC;
		 P0 : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT il_level1s
	PORT(LSZD_Pos0 : IN STD_LOGIC;
		 LSZD_Pos1 : IN STD_LOGIC;
		 Cout_0 : IN STD_LOGIC;
		 In_0 : IN STD_LOGIC;
		 In_1 : IN STD_LOGIC;
		 In_2 : IN STD_LOGIC;
		 pn1 : OUT STD_LOGIC;
		 Out_0 : OUT STD_LOGIC;
		 Out_1 : OUT STD_LOGIC;
		 Out_2 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lszd_level3
	PORT(MS0 : IN STD_LOGIC;
		 MS1 : IN STD_LOGIC;
		 MS2 : IN STD_LOGIC;
		 MSH_LSsumbit_2 : IN STD_LOGIC;
		 MSH_LSsumbit_1 : IN STD_LOGIC;
		 MSH_LSsumbit_0 : IN STD_LOGIC;
		 NZ_MS : IN STD_LOGIC;
		 NZ_LS : IN STD_LOGIC;
		 P3 : OUT STD_LOGIC;
		 P2 : OUT STD_LOGIC;
		 P1 : OUT STD_LOGIC;
		 P0 : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT il_level4_new
	PORT(LSZD_Pos0 : IN STD_LOGIC;
		 LSZD_Pos1 : IN STD_LOGIC;
		 LSZD_Pos2 : IN STD_LOGIC;
		 LSZD_Pos3 : IN STD_LOGIC;
		 LSZD_Pos4 : IN STD_LOGIC;
		 Cout_0 : IN STD_LOGIC;
		 In_0 : IN STD_LOGIC;
		 In_1 : IN STD_LOGIC;
		 In_2 : IN STD_LOGIC;
		 In_3 : IN STD_LOGIC;
		 In_4 : IN STD_LOGIC;
		 In_5 : IN STD_LOGIC;
		 In_6 : IN STD_LOGIC;
		 In_7 : IN STD_LOGIC;
		 In_8 : IN STD_LOGIC;
		 In_9 : IN STD_LOGIC;
		 In_10 : IN STD_LOGIC;
		 In_11 : IN STD_LOGIC;
		 In_12 : IN STD_LOGIC;
		 In_13 : IN STD_LOGIC;
		 In_14 : IN STD_LOGIC;
		 In_15 : IN STD_LOGIC;
		 In_16 : IN STD_LOGIC;
		 Out_0 : OUT STD_LOGIC;
		 Out_1 : OUT STD_LOGIC;
		 Out_2 : OUT STD_LOGIC;
		 Out_3 : OUT STD_LOGIC;
		 Out_4 : OUT STD_LOGIC;
		 Out_5 : OUT STD_LOGIC;
		 Out_6 : OUT STD_LOGIC;
		 Out_7 : OUT STD_LOGIC;
		 Out_8 : OUT STD_LOGIC;
		 Out_9 : OUT STD_LOGIC;
		 Out_10 : OUT STD_LOGIC;
		 Out_11 : OUT STD_LOGIC;
		 Out_12 : OUT STD_LOGIC;
		 Out_13 : OUT STD_LOGIC;
		 Out_14 : OUT STD_LOGIC;
		 Out_15 : OUT STD_LOGIC;
		 Out_16 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT il_level3_new
	PORT(LSZD_Pos0 : IN STD_LOGIC;
		 LSZD_Pos1 : IN STD_LOGIC;
		 LSZD_Pos2 : IN STD_LOGIC;
		 LSZD_Pos3 : IN STD_LOGIC;
		 NZFlag : IN STD_LOGIC;
		 Cout_0 : IN STD_LOGIC;
		 In_0 : IN STD_LOGIC;
		 In_1 : IN STD_LOGIC;
		 In_2 : IN STD_LOGIC;
		 In_3 : IN STD_LOGIC;
		 In_4 : IN STD_LOGIC;
		 In_5 : IN STD_LOGIC;
		 In_6 : IN STD_LOGIC;
		 In_7 : IN STD_LOGIC;
		 In_8 : IN STD_LOGIC;
		 Out_0 : OUT STD_LOGIC;
		 Out_1 : OUT STD_LOGIC;
		 Out_2 : OUT STD_LOGIC;
		 Out_3 : OUT STD_LOGIC;
		 Out_4 : OUT STD_LOGIC;
		 Out_5 : OUT STD_LOGIC;
		 Out_6 : OUT STD_LOGIC;
		 Out_7 : OUT STD_LOGIC;
		 Out_8 : OUT STD_LOGIC;
		 Out_9 : OUT STD_LOGIC;
		 Out_10 : OUT STD_LOGIC;
		 Out_11 : OUT STD_LOGIC;
		 Out_12 : OUT STD_LOGIC;
		 Out_13 : OUT STD_LOGIC;
		 Out_14 : OUT STD_LOGIC;
		 Out_15 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lszd_level4
	PORT(MS0 : IN STD_LOGIC;
		 MS1 : IN STD_LOGIC;
		 MS2 : IN STD_LOGIC;
		 MS3 : IN STD_LOGIC;
		 NZ_MS : IN STD_LOGIC;
		 NZ_LS : IN STD_LOGIC;
		 MSH_LSsumbit_0 : IN STD_LOGIC;
		 MSH_LSsumbit_1 : IN STD_LOGIC;
		 MSH_LSsumbit_2 : IN STD_LOGIC;
		 MSH_LSsumbit_3 : IN STD_LOGIC;
		 P4 : OUT STD_LOGIC;
		 P3 : OUT STD_LOGIC;
		 P2 : OUT STD_LOGIC;
		 P1 : OUT STD_LOGIC;
		 P0 : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lszd_level5
	PORT(MS0 : IN STD_LOGIC;
		 MS1 : IN STD_LOGIC;
		 MS2 : IN STD_LOGIC;
		 MS3 : IN STD_LOGIC;
		 MS4 : IN STD_LOGIC;
		 NZ_MS : IN STD_LOGIC;
		 NZ_LS : IN STD_LOGIC;
		 MSH_LSsumbit_0 : IN STD_LOGIC;
		 MSH_LSsumbit_1 : IN STD_LOGIC;
		 MSH_LSsumbit_2 : IN STD_LOGIC;
		 MSH_LSsumbit_3 : IN STD_LOGIC;
		 P5 : OUT STD_LOGIC;
		 P4 : OUT STD_LOGIC;
		 P3 : OUT STD_LOGIC;
		 P2 : OUT STD_LOGIC;
		 P1 : OUT STD_LOGIC;
		 P0 : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lszd_level2_new
	PORT(MS0 : IN STD_LOGIC;
		 MS1 : IN STD_LOGIC;
		 MSH_LSsumbit_1 : IN STD_LOGIC;
		 MSH_LSsumbit_0 : IN STD_LOGIC;
		 NZ_MS : IN STD_LOGIC;
		 NZ_LS : IN STD_LOGIC;
		 P2 : OUT STD_LOGIC;
		 P1 : OUT STD_LOGIC;
		 P0 : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT leaf_cin
	PORT(A_1 : IN STD_LOGIC;
		 B_1 : IN STD_LOGIC;
		 A_0 : IN STD_LOGIC;
		 B_0 : IN STD_LOGIC;
		 Cin_init : IN STD_LOGIC;
		 Sum_1p : OUT STD_LOGIC;
		 Cout_1p : OUT STD_LOGIC;
		 NZ : OUT STD_LOGIC;
		 Sum_0 : OUT STD_LOGIC;
		 Pos : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	sum_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(64 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_490 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_491 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_492 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_493 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_494 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_495 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_496 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_497 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_498 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_499 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_500 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_501 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_502 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_503 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_504 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_505 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_506 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_507 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_508 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_509 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_510 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_511 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_512 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_513 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_514 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_515 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_516 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_517 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_518 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_519 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_520 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_521 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_522 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_523 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_524 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_525 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_526 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_527 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_528 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_529 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_530 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_531 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_532 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_533 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_534 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_535 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_178 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_182 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_183 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_184 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_185 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_186 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_187 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_198 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_202 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_203 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_204 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_205 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_536 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_207 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_537 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_538 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_539 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_212 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_213 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_214 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_215 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_216 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_540 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_220 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_541 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_224 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_225 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_228 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_229 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_542 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_232 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_233 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_236 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_543 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_240 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_247 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_248 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_249 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_250 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_251 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_252 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_544 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_545 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_255 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_256 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_546 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_547 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_260 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_548 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_262 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_264 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_549 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_266 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_267 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_268 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_270 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_271 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_550 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_551 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_552 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_278 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_279 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_280 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_281 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_282 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_553 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_554 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_555 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_556 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_289 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_557 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_558 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_292 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_293 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_294 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_295 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_297 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_298 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_299 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_559 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_301 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_302 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_560 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_561 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_562 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_563 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_564 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_308 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_565 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_566 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_567 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_312 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_313 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_314 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_315 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_316 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_317 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_324 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_325 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_568 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_569 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_570 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_571 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_572 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_331 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_573 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_574 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_575 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_576 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_336 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_337 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_338 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_339 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_340 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_341 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_342 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_343 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_344 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_345 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_346 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_347 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_348 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_359 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_360 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_361 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_362 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_577 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_578 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_365 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_366 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_367 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_373 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_374 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_579 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_580 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_383 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_384 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_581 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_582 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_583 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_584 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_389 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_390 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_395 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_396 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_400 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_403 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_404 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_405 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_585 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_586 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_410 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_411 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_416 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_417 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_587 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_588 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_422 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_423 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_428 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_429 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_589 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_590 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_434 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_435 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_438 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_440 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_441 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_442 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_443 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_444 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_446 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_447 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_448 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_449 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_450 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_452 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_453 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_456 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_458 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_459 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_460 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_461 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_462 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_464 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_465 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_468 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_470 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_471 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_472 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_473 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_474 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_476 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_477 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_480 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_482 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_483 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_486 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_488 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_489 :  STD_LOGIC;


BEGIN 



b2v_inst : il_level5_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_0,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_1,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_2,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_3,
		 LSZD_Pos4 => SYNTHESIZED_WIRE_4,
		 LSZD_Pos5 => SYNTHESIZED_WIRE_5,
		 NZFlag => SYNTHESIZED_WIRE_6,
		 Cout_0 => SYNTHESIZED_WIRE_7,
		 In_0 => SYNTHESIZED_WIRE_490,
		 In_1 => SYNTHESIZED_WIRE_491,
		 In_2 => SYNTHESIZED_WIRE_492,
		 In_3 => SYNTHESIZED_WIRE_493,
		 In_4 => SYNTHESIZED_WIRE_12,
		 In_5 => SYNTHESIZED_WIRE_13,
		 In_6 => SYNTHESIZED_WIRE_14,
		 In_7 => SYNTHESIZED_WIRE_15,
		 In_8 => SYNTHESIZED_WIRE_16,
		 In_9 => SYNTHESIZED_WIRE_17,
		 In_10 => SYNTHESIZED_WIRE_18,
		 In_11 => SYNTHESIZED_WIRE_19,
		 In_12 => SYNTHESIZED_WIRE_20,
		 In_13 => SYNTHESIZED_WIRE_21,
		 In_14 => SYNTHESIZED_WIRE_22,
		 In_15 => SYNTHESIZED_WIRE_23,
		 In_16 => SYNTHESIZED_WIRE_24,
		 In_17 => SYNTHESIZED_WIRE_25,
		 In_18 => SYNTHESIZED_WIRE_26,
		 In_19 => SYNTHESIZED_WIRE_27,
		 In_20 => SYNTHESIZED_WIRE_28,
		 In_21 => SYNTHESIZED_WIRE_29,
		 In_22 => SYNTHESIZED_WIRE_30,
		 In_23 => SYNTHESIZED_WIRE_31,
		 In_24 => SYNTHESIZED_WIRE_32,
		 In_25 => SYNTHESIZED_WIRE_33,
		 In_26 => SYNTHESIZED_WIRE_34,
		 In_27 => SYNTHESIZED_WIRE_35,
		 In_28 => SYNTHESIZED_WIRE_36,
		 In_29 => SYNTHESIZED_WIRE_37,
		 In_30 => SYNTHESIZED_WIRE_38,
		 In_31 => SYNTHESIZED_WIRE_39,
		 In_32 => SYNTHESIZED_WIRE_40,
		 Out_0 => sum_ALTERA_SYNTHESIZED(32),
		 Out_1 => sum_ALTERA_SYNTHESIZED(33),
		 Out_2 => sum_ALTERA_SYNTHESIZED(34),
		 Out_3 => sum_ALTERA_SYNTHESIZED(35),
		 Out_4 => sum_ALTERA_SYNTHESIZED(36),
		 Out_5 => sum_ALTERA_SYNTHESIZED(37),
		 Out_6 => sum_ALTERA_SYNTHESIZED(38),
		 Out_7 => sum_ALTERA_SYNTHESIZED(39),
		 Out_8 => sum_ALTERA_SYNTHESIZED(40),
		 Out_9 => sum_ALTERA_SYNTHESIZED(41),
		 Out_10 => sum_ALTERA_SYNTHESIZED(42),
		 Out_11 => sum_ALTERA_SYNTHESIZED(43),
		 Out_12 => sum_ALTERA_SYNTHESIZED(44),
		 Out_13 => sum_ALTERA_SYNTHESIZED(45),
		 Out_14 => sum_ALTERA_SYNTHESIZED(46),
		 Out_15 => sum_ALTERA_SYNTHESIZED(47),
		 Out_16 => sum_ALTERA_SYNTHESIZED(48),
		 Out_17 => sum_ALTERA_SYNTHESIZED(49),
		 Out_18 => sum_ALTERA_SYNTHESIZED(50),
		 Out_19 => sum_ALTERA_SYNTHESIZED(51),
		 Out_20 => sum_ALTERA_SYNTHESIZED(52),
		 Out_21 => sum_ALTERA_SYNTHESIZED(53),
		 Out_22 => sum_ALTERA_SYNTHESIZED(54),
		 Out_23 => sum_ALTERA_SYNTHESIZED(55),
		 Out_24 => sum_ALTERA_SYNTHESIZED(56),
		 Out_25 => sum_ALTERA_SYNTHESIZED(57),
		 Out_26 => sum_ALTERA_SYNTHESIZED(58),
		 Out_27 => sum_ALTERA_SYNTHESIZED(59),
		 Out_28 => sum_ALTERA_SYNTHESIZED(60),
		 Out_29 => sum_ALTERA_SYNTHESIZED(61),
		 Out_30 => sum_ALTERA_SYNTHESIZED(62),
		 Out_31 => sum_ALTERA_SYNTHESIZED(63),
		 Out_32 => sum_ALTERA_SYNTHESIZED(64));


b2v_inst1 : leaf
PORT MAP(A_1 => a(43),
		 B_1 => b(43),
		 A_0 => a(42),
		 B_0 => b(42),
		 Sum_1p => SYNTHESIZED_WIRE_118,
		 Cout_1p => SYNTHESIZED_WIRE_119,
		 NZ => SYNTHESIZED_WIRE_200,
		 Sum_0 => SYNTHESIZED_WIRE_517,
		 Pos => SYNTHESIZED_WIRE_198);


b2v_inst10 : leaf
PORT MAP(A_1 => a(13),
		 B_1 => b(13),
		 A_0 => a(12),
		 B_0 => b(12),
		 Sum_1p => SYNTHESIZED_WIRE_583,
		 Cout_1p => SYNTHESIZED_WIRE_438,
		 NZ => SYNTHESIZED_WIRE_224,
		 Sum_0 => SYNTHESIZED_WIRE_584);


b2v_inst11 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_41,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_42,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_43,
		 Cout_0 => SYNTHESIZED_WIRE_44,
		 In_0 => SYNTHESIZED_WIRE_494,
		 In_1 => SYNTHESIZED_WIRE_495,
		 In_2 => SYNTHESIZED_WIRE_47,
		 In_3 => SYNTHESIZED_WIRE_48,
		 In_4 => SYNTHESIZED_WIRE_49,
		 Out_0 => SYNTHESIZED_WIRE_142,
		 Out_1 => SYNTHESIZED_WIRE_141,
		 Out_2 => SYNTHESIZED_WIRE_140,
		 Out_3 => SYNTHESIZED_WIRE_139,
		 Out_4 => SYNTHESIZED_WIRE_178);


b2v_inst12 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_50,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_496,
		 NZ_MS => SYNTHESIZED_WIRE_52,
		 NZ_LS => SYNTHESIZED_WIRE_53,
		 P1 => SYNTHESIZED_WIRE_443,
		 P0 => SYNTHESIZED_WIRE_442,
		 NZ => SYNTHESIZED_WIRE_384);


b2v_inst13 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_54,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_497,
		 NZ_MS => SYNTHESIZED_WIRE_56,
		 NZ_LS => SYNTHESIZED_WIRE_57,
		 P1 => SYNTHESIZED_WIRE_153,
		 P0 => SYNTHESIZED_WIRE_152,
		 NZ => SYNTHESIZED_WIRE_390);


b2v_inst14 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_498,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_499,
		 Cout_0 => SYNTHESIZED_WIRE_60,
		 In_0 => SYNTHESIZED_WIRE_500,
		 In_1 => SYNTHESIZED_WIRE_62,
		 In_2 => SYNTHESIZED_WIRE_63,
		 Out_0 => SYNTHESIZED_WIRE_47,
		 Out_1 => SYNTHESIZED_WIRE_48,
		 Out_2 => SYNTHESIZED_WIRE_49);


b2v_inst15 : leaf
PORT MAP(A_1 => a(23),
		 B_1 => b(23),
		 A_0 => a(22),
		 B_0 => b(22),
		 Sum_1p => SYNTHESIZED_WIRE_62,
		 Cout_1p => SYNTHESIZED_WIRE_63,
		 NZ => SYNTHESIZED_WIRE_227,
		 Sum_0 => SYNTHESIZED_WIRE_500,
		 Pos => SYNTHESIZED_WIRE_225);


b2v_inst16 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_64,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_501,
		 NZ_MS => SYNTHESIZED_WIRE_66,
		 NZ_LS => SYNTHESIZED_WIRE_67,
		 P1 => SYNTHESIZED_WIRE_449,
		 P0 => SYNTHESIZED_WIRE_448,
		 NZ => SYNTHESIZED_WIRE_396);


b2v_inst17 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_68,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_69,
		 Cout_0 => SYNTHESIZED_WIRE_70,
		 In_0 => SYNTHESIZED_WIRE_502,
		 In_1 => SYNTHESIZED_WIRE_72,
		 In_2 => SYNTHESIZED_WIRE_73,
		 Out_0 => SYNTHESIZED_WIRE_508,
		 Out_1 => SYNTHESIZED_WIRE_182,
		 Out_2 => SYNTHESIZED_WIRE_77);


b2v_inst18 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_503,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_504,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_505,
		 Cout_0 => SYNTHESIZED_WIRE_77,
		 In_0 => SYNTHESIZED_WIRE_506,
		 In_1 => SYNTHESIZED_WIRE_507,
		 In_2 => SYNTHESIZED_WIRE_80,
		 In_3 => SYNTHESIZED_WIRE_81,
		 In_4 => SYNTHESIZED_WIRE_82,
		 Out_0 => SYNTHESIZED_WIRE_183,
		 Out_1 => SYNTHESIZED_WIRE_184,
		 Out_2 => SYNTHESIZED_WIRE_185,
		 Out_3 => SYNTHESIZED_WIRE_186,
		 Out_4 => SYNTHESIZED_WIRE_187);


b2v_inst19 : leaf
PORT MAP(A_1 => a(29),
		 B_1 => b(29),
		 A_0 => a(28),
		 B_0 => b(28),
		 Sum_1p => SYNTHESIZED_WIRE_507,
		 Cout_1p => SYNTHESIZED_WIRE_456,
		 NZ => SYNTHESIZED_WIRE_232,
		 Sum_0 => SYNTHESIZED_WIRE_506);


b2v_inst2 : leaf
PORT MAP(A_1 => a(9),
		 B_1 => b(9),
		 A_0 => a(8),
		 B_0 => b(8),
		 Sum_1p => SYNTHESIZED_WIRE_529,
		 Cout_1p => SYNTHESIZED_WIRE_154,
		 NZ => SYNTHESIZED_WIRE_57,
		 Sum_0 => SYNTHESIZED_WIRE_528);


b2v_inst20 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_83,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_502,
		 NZ_MS => SYNTHESIZED_WIRE_85,
		 NZ_LS => SYNTHESIZED_WIRE_86,
		 P1 => SYNTHESIZED_WIRE_69,
		 P0 => SYNTHESIZED_WIRE_68,
		 NZ => SYNTHESIZED_WIRE_411);


b2v_inst21 : leaf
PORT MAP(A_1 => a(25),
		 B_1 => b(25),
		 A_0 => a(24),
		 B_0 => b(24),
		 Sum_1p => SYNTHESIZED_WIRE_509,
		 Cout_1p => SYNTHESIZED_WIRE_70,
		 NZ => SYNTHESIZED_WIRE_86,
		 Sum_0 => SYNTHESIZED_WIRE_510);


b2v_inst22 : lszd_level3
PORT MAP(MS0 => SYNTHESIZED_WIRE_503,
		 MS1 => SYNTHESIZED_WIRE_504,
		 MS2 => SYNTHESIZED_WIRE_505,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_508,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_509,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_510,
		 NZ_MS => SYNTHESIZED_WIRE_93,
		 NZ_LS => SYNTHESIZED_WIRE_94,
		 P3 => SYNTHESIZED_WIRE_534,
		 P2 => SYNTHESIZED_WIRE_533,
		 P1 => SYNTHESIZED_WIRE_532,
		 P0 => SYNTHESIZED_WIRE_531,
		 NZ => SYNTHESIZED_WIRE_535);


b2v_inst23 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_95,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_96,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_97,
		 Cout_0 => SYNTHESIZED_WIRE_98,
		 In_0 => SYNTHESIZED_WIRE_511,
		 In_1 => SYNTHESIZED_WIRE_512,
		 In_2 => SYNTHESIZED_WIRE_101,
		 In_3 => SYNTHESIZED_WIRE_102,
		 In_4 => SYNTHESIZED_WIRE_103,
		 Out_0 => SYNTHESIZED_WIRE_15,
		 Out_1 => SYNTHESIZED_WIRE_14,
		 Out_2 => SYNTHESIZED_WIRE_13,
		 Out_3 => SYNTHESIZED_WIRE_12,
		 Out_4 => SYNTHESIZED_WIRE_207);


b2v_inst24 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_513,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_514,
		 Cout_0 => SYNTHESIZED_WIRE_106,
		 In_0 => SYNTHESIZED_WIRE_515,
		 In_1 => SYNTHESIZED_WIRE_108,
		 In_2 => SYNTHESIZED_WIRE_109,
		 Out_0 => SYNTHESIZED_WIRE_101,
		 Out_1 => SYNTHESIZED_WIRE_102,
		 Out_2 => SYNTHESIZED_WIRE_103);


b2v_inst25 : leaf
PORT MAP(A_1 => a(39),
		 B_1 => b(39),
		 A_0 => a(38),
		 B_0 => b(38),
		 Sum_1p => SYNTHESIZED_WIRE_108,
		 Cout_1p => SYNTHESIZED_WIRE_109,
		 NZ => SYNTHESIZED_WIRE_235,
		 Sum_0 => SYNTHESIZED_WIRE_515,
		 Pos => SYNTHESIZED_WIRE_233);


b2v_inst26 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_110,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_516,
		 NZ_MS => SYNTHESIZED_WIRE_112,
		 NZ_LS => SYNTHESIZED_WIRE_113,
		 P1 => SYNTHESIZED_WIRE_461,
		 P0 => SYNTHESIZED_WIRE_460,
		 NZ => SYNTHESIZED_WIRE_417);


b2v_inst27 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_114,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_115,
		 Cout_0 => SYNTHESIZED_WIRE_116,
		 In_0 => SYNTHESIZED_WIRE_517,
		 In_1 => SYNTHESIZED_WIRE_118,
		 In_2 => SYNTHESIZED_WIRE_119,
		 Out_0 => SYNTHESIZED_WIRE_539,
		 Out_1 => SYNTHESIZED_WIRE_211,
		 Out_2 => SYNTHESIZED_WIRE_123);


b2v_inst28 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_518,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_519,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_520,
		 Cout_0 => SYNTHESIZED_WIRE_123,
		 In_0 => SYNTHESIZED_WIRE_521,
		 In_1 => SYNTHESIZED_WIRE_522,
		 In_2 => SYNTHESIZED_WIRE_126,
		 In_3 => SYNTHESIZED_WIRE_127,
		 In_4 => SYNTHESIZED_WIRE_128,
		 Out_0 => SYNTHESIZED_WIRE_212,
		 Out_1 => SYNTHESIZED_WIRE_213,
		 Out_2 => SYNTHESIZED_WIRE_214,
		 Out_3 => SYNTHESIZED_WIRE_215,
		 Out_4 => SYNTHESIZED_WIRE_216);


b2v_inst29 : il_level4_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_129,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_130,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_131,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_132,
		 LSZD_Pos4 => SYNTHESIZED_WIRE_133,
		 Cout_0 => SYNTHESIZED_WIRE_134,
		 In_0 => SYNTHESIZED_WIRE_523,
		 In_1 => SYNTHESIZED_WIRE_524,
		 In_2 => SYNTHESIZED_WIRE_525,
		 In_3 => SYNTHESIZED_WIRE_526,
		 In_4 => SYNTHESIZED_WIRE_139,
		 In_5 => SYNTHESIZED_WIRE_140,
		 In_6 => SYNTHESIZED_WIRE_141,
		 In_7 => SYNTHESIZED_WIRE_142,
		 In_8 => SYNTHESIZED_WIRE_143,
		 In_9 => SYNTHESIZED_WIRE_144,
		 In_10 => SYNTHESIZED_WIRE_145,
		 In_11 => SYNTHESIZED_WIRE_146,
		 In_12 => SYNTHESIZED_WIRE_147,
		 In_13 => SYNTHESIZED_WIRE_148,
		 In_14 => SYNTHESIZED_WIRE_149,
		 In_15 => SYNTHESIZED_WIRE_150,
		 In_16 => SYNTHESIZED_WIRE_151,
		 Out_0 => sum_ALTERA_SYNTHESIZED(16),
		 Out_1 => sum_ALTERA_SYNTHESIZED(17),
		 Out_2 => sum_ALTERA_SYNTHESIZED(18),
		 Out_3 => sum_ALTERA_SYNTHESIZED(19),
		 Out_4 => sum_ALTERA_SYNTHESIZED(20),
		 Out_5 => sum_ALTERA_SYNTHESIZED(21),
		 Out_6 => sum_ALTERA_SYNTHESIZED(22),
		 Out_7 => sum_ALTERA_SYNTHESIZED(23),
		 Out_8 => sum_ALTERA_SYNTHESIZED(24),
		 Out_9 => sum_ALTERA_SYNTHESIZED(25),
		 Out_10 => sum_ALTERA_SYNTHESIZED(26),
		 Out_11 => sum_ALTERA_SYNTHESIZED(27),
		 Out_12 => sum_ALTERA_SYNTHESIZED(28),
		 Out_13 => sum_ALTERA_SYNTHESIZED(29),
		 Out_14 => sum_ALTERA_SYNTHESIZED(30),
		 Out_15 => sum_ALTERA_SYNTHESIZED(31),
		 Out_16 => SYNTHESIZED_WIRE_7);


b2v_inst3 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_152,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_153,
		 Cout_0 => SYNTHESIZED_WIRE_154,
		 In_0 => SYNTHESIZED_WIRE_497,
		 In_1 => SYNTHESIZED_WIRE_156,
		 In_2 => SYNTHESIZED_WIRE_157,
		 Out_0 => SYNTHESIZED_WIRE_530,
		 Out_1 => SYNTHESIZED_WIRE_167,
		 Out_2 => SYNTHESIZED_WIRE_400);


b2v_inst30 : il_level3_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_158,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_159,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_160,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_161,
		 NZFlag => SYNTHESIZED_WIRE_527,
		 Cout_0 => SYNTHESIZED_WIRE_163,
		 In_0 => SYNTHESIZED_WIRE_528,
		 In_1 => SYNTHESIZED_WIRE_529,
		 In_2 => SYNTHESIZED_WIRE_530,
		 In_3 => SYNTHESIZED_WIRE_167,
		 In_4 => SYNTHESIZED_WIRE_168,
		 In_5 => SYNTHESIZED_WIRE_169,
		 In_6 => SYNTHESIZED_WIRE_170,
		 In_7 => SYNTHESIZED_WIRE_171,
		 In_8 => SYNTHESIZED_WIRE_172,
		 Out_0 => sum_ALTERA_SYNTHESIZED(8),
		 Out_1 => sum_ALTERA_SYNTHESIZED(9),
		 Out_2 => sum_ALTERA_SYNTHESIZED(10),
		 Out_3 => sum_ALTERA_SYNTHESIZED(11),
		 Out_4 => sum_ALTERA_SYNTHESIZED(12),
		 Out_5 => sum_ALTERA_SYNTHESIZED(13),
		 Out_6 => sum_ALTERA_SYNTHESIZED(14),
		 Out_7 => sum_ALTERA_SYNTHESIZED(15),
		 Out_8 => SYNTHESIZED_WIRE_134);


b2v_inst31 : il_level3_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_531,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_532,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_533,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_534,
		 NZFlag => SYNTHESIZED_WIRE_535,
		 Cout_0 => SYNTHESIZED_WIRE_178,
		 In_0 => SYNTHESIZED_WIRE_510,
		 In_1 => SYNTHESIZED_WIRE_509,
		 In_2 => SYNTHESIZED_WIRE_508,
		 In_3 => SYNTHESIZED_WIRE_182,
		 In_4 => SYNTHESIZED_WIRE_183,
		 In_5 => SYNTHESIZED_WIRE_184,
		 In_6 => SYNTHESIZED_WIRE_185,
		 In_7 => SYNTHESIZED_WIRE_186,
		 In_8 => SYNTHESIZED_WIRE_187,
		 Out_0 => SYNTHESIZED_WIRE_143,
		 Out_1 => SYNTHESIZED_WIRE_144,
		 Out_2 => SYNTHESIZED_WIRE_145,
		 Out_3 => SYNTHESIZED_WIRE_146,
		 Out_4 => SYNTHESIZED_WIRE_147,
		 Out_5 => SYNTHESIZED_WIRE_148,
		 Out_6 => SYNTHESIZED_WIRE_149,
		 Out_7 => SYNTHESIZED_WIRE_150,
		 Out_8 => SYNTHESIZED_WIRE_151);


b2v_inst32 : lszd_level4
PORT MAP(MS0 => SYNTHESIZED_WIRE_531,
		 MS1 => SYNTHESIZED_WIRE_532,
		 MS2 => SYNTHESIZED_WIRE_533,
		 MS3 => SYNTHESIZED_WIRE_534,
		 NZ_MS => SYNTHESIZED_WIRE_535,
		 NZ_LS => SYNTHESIZED_WIRE_527,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_523,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_524,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_525,
		 MSH_LSsumbit_3 => SYNTHESIZED_WIRE_526,
		 P4 => SYNTHESIZED_WIRE_133,
		 P3 => SYNTHESIZED_WIRE_132,
		 P2 => SYNTHESIZED_WIRE_131,
		 P1 => SYNTHESIZED_WIRE_130,
		 P0 => SYNTHESIZED_WIRE_129,
		 NZ => SYNTHESIZED_WIRE_374);


b2v_inst33 : leaf
PORT MAP(A_1 => a(45),
		 B_1 => b(45),
		 A_0 => a(44),
		 B_0 => b(44),
		 Sum_1p => SYNTHESIZED_WIRE_522,
		 Cout_1p => SYNTHESIZED_WIRE_468,
		 NZ => SYNTHESIZED_WIRE_240,
		 Sum_0 => SYNTHESIZED_WIRE_521);


b2v_inst34 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_198,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_517,
		 NZ_MS => SYNTHESIZED_WIRE_200,
		 NZ_LS => SYNTHESIZED_WIRE_201,
		 P1 => SYNTHESIZED_WIRE_115,
		 P0 => SYNTHESIZED_WIRE_114,
		 NZ => SYNTHESIZED_WIRE_423);


b2v_inst35 : leaf
PORT MAP(A_1 => a(41),
		 B_1 => b(41),
		 A_0 => a(40),
		 B_0 => b(40),
		 Sum_1p => SYNTHESIZED_WIRE_538,
		 Cout_1p => SYNTHESIZED_WIRE_116,
		 NZ => SYNTHESIZED_WIRE_201,
		 Sum_0 => SYNTHESIZED_WIRE_537);


b2v_inst36 : il_level3_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_202,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_203,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_204,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_205,
		 NZFlag => SYNTHESIZED_WIRE_536,
		 Cout_0 => SYNTHESIZED_WIRE_207,
		 In_0 => SYNTHESIZED_WIRE_537,
		 In_1 => SYNTHESIZED_WIRE_538,
		 In_2 => SYNTHESIZED_WIRE_539,
		 In_3 => SYNTHESIZED_WIRE_211,
		 In_4 => SYNTHESIZED_WIRE_212,
		 In_5 => SYNTHESIZED_WIRE_213,
		 In_6 => SYNTHESIZED_WIRE_214,
		 In_7 => SYNTHESIZED_WIRE_215,
		 In_8 => SYNTHESIZED_WIRE_216,
		 Out_0 => SYNTHESIZED_WIRE_23,
		 Out_1 => SYNTHESIZED_WIRE_22,
		 Out_2 => SYNTHESIZED_WIRE_21,
		 Out_3 => SYNTHESIZED_WIRE_20,
		 Out_4 => SYNTHESIZED_WIRE_19,
		 Out_5 => SYNTHESIZED_WIRE_18,
		 Out_6 => SYNTHESIZED_WIRE_17,
		 Out_7 => SYNTHESIZED_WIRE_16,
		 Out_8 => SYNTHESIZED_WIRE_331);


b2v_inst37 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_217,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_540,
		 NZ_MS => SYNTHESIZED_WIRE_219,
		 NZ_LS => SYNTHESIZED_WIRE_220,
		 P1 => SYNTHESIZED_WIRE_580,
		 P0 => SYNTHESIZED_WIRE_579,
		 NZ => SYNTHESIZED_WIRE_383);


b2v_inst38 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_221,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_541,
		 NZ_MS => SYNTHESIZED_WIRE_223,
		 NZ_LS => SYNTHESIZED_WIRE_224,
		 P1 => SYNTHESIZED_WIRE_582,
		 P0 => SYNTHESIZED_WIRE_581,
		 NZ => SYNTHESIZED_WIRE_389);


b2v_inst39 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_225,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_500,
		 NZ_MS => SYNTHESIZED_WIRE_227,
		 NZ_LS => SYNTHESIZED_WIRE_228,
		 P1 => SYNTHESIZED_WIRE_499,
		 P0 => SYNTHESIZED_WIRE_498,
		 NZ => SYNTHESIZED_WIRE_395);


b2v_inst4 : leaf
PORT MAP(A_1 => a(27),
		 B_1 => b(27),
		 A_0 => a(26),
		 B_0 => b(26),
		 Sum_1p => SYNTHESIZED_WIRE_72,
		 Cout_1p => SYNTHESIZED_WIRE_73,
		 NZ => SYNTHESIZED_WIRE_85,
		 Sum_0 => SYNTHESIZED_WIRE_502,
		 Pos => SYNTHESIZED_WIRE_83);


b2v_inst40 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_229,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_542,
		 NZ_MS => SYNTHESIZED_WIRE_231,
		 NZ_LS => SYNTHESIZED_WIRE_232,
		 P1 => SYNTHESIZED_WIRE_586,
		 P0 => SYNTHESIZED_WIRE_585,
		 NZ => SYNTHESIZED_WIRE_410);


b2v_inst41 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_233,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_515,
		 NZ_MS => SYNTHESIZED_WIRE_235,
		 NZ_LS => SYNTHESIZED_WIRE_236,
		 P1 => SYNTHESIZED_WIRE_514,
		 P0 => SYNTHESIZED_WIRE_513,
		 NZ => SYNTHESIZED_WIRE_416);


b2v_inst42 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_237,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_543,
		 NZ_MS => SYNTHESIZED_WIRE_239,
		 NZ_LS => SYNTHESIZED_WIRE_240,
		 P1 => SYNTHESIZED_WIRE_588,
		 P0 => SYNTHESIZED_WIRE_587,
		 NZ => SYNTHESIZED_WIRE_422);


b2v_inst43 : lszd_level3
PORT MAP(MS0 => SYNTHESIZED_WIRE_518,
		 MS1 => SYNTHESIZED_WIRE_519,
		 MS2 => SYNTHESIZED_WIRE_520,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_539,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_538,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_537,
		 NZ_MS => SYNTHESIZED_WIRE_247,
		 NZ_LS => SYNTHESIZED_WIRE_248,
		 P3 => SYNTHESIZED_WIRE_205,
		 P2 => SYNTHESIZED_WIRE_204,
		 P1 => SYNTHESIZED_WIRE_203,
		 P0 => SYNTHESIZED_WIRE_202,
		 NZ => SYNTHESIZED_WIRE_536);


b2v_inst44 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_249,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_250,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_251,
		 Cout_0 => SYNTHESIZED_WIRE_252,
		 In_0 => SYNTHESIZED_WIRE_544,
		 In_1 => SYNTHESIZED_WIRE_545,
		 In_2 => SYNTHESIZED_WIRE_255,
		 In_3 => SYNTHESIZED_WIRE_256,
		 In_4 => SYNTHESIZED_WIRE_257,
		 Out_0 => SYNTHESIZED_WIRE_339,
		 Out_1 => SYNTHESIZED_WIRE_338,
		 Out_2 => SYNTHESIZED_WIRE_337,
		 Out_3 => SYNTHESIZED_WIRE_336,
		 Out_4 => SYNTHESIZED_WIRE_308);


b2v_inst45 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_546,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_547,
		 Cout_0 => SYNTHESIZED_WIRE_260,
		 In_0 => SYNTHESIZED_WIRE_548,
		 In_1 => SYNTHESIZED_WIRE_262,
		 In_2 => SYNTHESIZED_WIRE_263,
		 Out_0 => SYNTHESIZED_WIRE_255,
		 Out_1 => SYNTHESIZED_WIRE_256,
		 Out_2 => SYNTHESIZED_WIRE_257);


b2v_inst46 : leaf
PORT MAP(A_1 => a(55),
		 B_1 => b(55),
		 A_0 => a(54),
		 B_0 => b(54),
		 Sum_1p => SYNTHESIZED_WIRE_262,
		 Cout_1p => SYNTHESIZED_WIRE_263,
		 NZ => SYNTHESIZED_WIRE_270,
		 Sum_0 => SYNTHESIZED_WIRE_548,
		 Pos => SYNTHESIZED_WIRE_268);


b2v_inst47 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_264,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_549,
		 NZ_MS => SYNTHESIZED_WIRE_266,
		 NZ_LS => SYNTHESIZED_WIRE_267,
		 P1 => SYNTHESIZED_WIRE_473,
		 P0 => SYNTHESIZED_WIRE_472,
		 NZ => SYNTHESIZED_WIRE_429);


b2v_inst48 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_268,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_548,
		 NZ_MS => SYNTHESIZED_WIRE_270,
		 NZ_LS => SYNTHESIZED_WIRE_271,
		 P1 => SYNTHESIZED_WIRE_547,
		 P0 => SYNTHESIZED_WIRE_546,
		 NZ => SYNTHESIZED_WIRE_428);


b2v_inst49 : leaf
PORT MAP(A_1 => a(59),
		 B_1 => b(59),
		 A_0 => a(58),
		 B_0 => b(58),
		 Sum_1p => SYNTHESIZED_WIRE_284,
		 Cout_1p => SYNTHESIZED_WIRE_285,
		 NZ => SYNTHESIZED_WIRE_297,
		 Sum_0 => SYNTHESIZED_WIRE_553,
		 Pos => SYNTHESIZED_WIRE_295);


b2v_inst5 : lszd_level3
PORT MAP(MS0 => SYNTHESIZED_WIRE_550,
		 MS1 => SYNTHESIZED_WIRE_551,
		 MS2 => SYNTHESIZED_WIRE_552,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_530,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_529,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_528,
		 NZ_MS => SYNTHESIZED_WIRE_278,
		 NZ_LS => SYNTHESIZED_WIRE_279,
		 P3 => SYNTHESIZED_WIRE_161,
		 P2 => SYNTHESIZED_WIRE_160,
		 P1 => SYNTHESIZED_WIRE_159,
		 P0 => SYNTHESIZED_WIRE_158,
		 NZ => SYNTHESIZED_WIRE_527);


b2v_inst50 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_280,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_281,
		 Cout_0 => SYNTHESIZED_WIRE_282,
		 In_0 => SYNTHESIZED_WIRE_553,
		 In_1 => SYNTHESIZED_WIRE_284,
		 In_2 => SYNTHESIZED_WIRE_285,
		 Out_0 => SYNTHESIZED_WIRE_567,
		 Out_1 => SYNTHESIZED_WIRE_312,
		 Out_2 => SYNTHESIZED_WIRE_289);


b2v_inst51 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_554,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_555,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_556,
		 Cout_0 => SYNTHESIZED_WIRE_289,
		 In_0 => SYNTHESIZED_WIRE_557,
		 In_1 => SYNTHESIZED_WIRE_558,
		 In_2 => SYNTHESIZED_WIRE_292,
		 In_3 => SYNTHESIZED_WIRE_293,
		 In_4 => SYNTHESIZED_WIRE_294,
		 Out_0 => SYNTHESIZED_WIRE_313,
		 Out_1 => SYNTHESIZED_WIRE_314,
		 Out_2 => SYNTHESIZED_WIRE_315,
		 Out_3 => SYNTHESIZED_WIRE_316,
		 Out_4 => SYNTHESIZED_WIRE_317);


b2v_inst52 : leaf
PORT MAP(A_1 => a(61),
		 B_1 => b(61),
		 A_0 => a(60),
		 B_0 => b(60),
		 Sum_1p => SYNTHESIZED_WIRE_558,
		 Cout_1p => SYNTHESIZED_WIRE_480,
		 NZ => SYNTHESIZED_WIRE_302,
		 Sum_0 => SYNTHESIZED_WIRE_557);


b2v_inst53 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_295,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_553,
		 NZ_MS => SYNTHESIZED_WIRE_297,
		 NZ_LS => SYNTHESIZED_WIRE_298,
		 P1 => SYNTHESIZED_WIRE_281,
		 P0 => SYNTHESIZED_WIRE_280,
		 NZ => SYNTHESIZED_WIRE_435);


b2v_inst54 : lszd_level1
PORT MAP(MS0 => SYNTHESIZED_WIRE_299,
		 MSH_LS_sumbit => SYNTHESIZED_WIRE_559,
		 NZ_MS => SYNTHESIZED_WIRE_301,
		 NZ_LS => SYNTHESIZED_WIRE_302,
		 P1 => SYNTHESIZED_WIRE_590,
		 P0 => SYNTHESIZED_WIRE_589,
		 NZ => SYNTHESIZED_WIRE_434);


b2v_inst55 : leaf
PORT MAP(A_1 => a(57),
		 B_1 => b(57),
		 A_0 => a(56),
		 B_0 => b(56),
		 Sum_1p => SYNTHESIZED_WIRE_566,
		 Cout_1p => SYNTHESIZED_WIRE_282,
		 NZ => SYNTHESIZED_WIRE_298,
		 Sum_0 => SYNTHESIZED_WIRE_565);


b2v_inst555 : leaf
PORT MAP(A_1 => a(11),
		 B_1 => b(11),
		 A_0 => a(10),
		 B_0 => b(10),
		 Sum_1p => SYNTHESIZED_WIRE_156,
		 Cout_1p => SYNTHESIZED_WIRE_157,
		 NZ => SYNTHESIZED_WIRE_56,
		 Sum_0 => SYNTHESIZED_WIRE_497,
		 Pos => SYNTHESIZED_WIRE_54);


b2v_inst56 : il_level3_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_560,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_561,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_562,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_563,
		 NZFlag => SYNTHESIZED_WIRE_564,
		 Cout_0 => SYNTHESIZED_WIRE_308,
		 In_0 => SYNTHESIZED_WIRE_565,
		 In_1 => SYNTHESIZED_WIRE_566,
		 In_2 => SYNTHESIZED_WIRE_567,
		 In_3 => SYNTHESIZED_WIRE_312,
		 In_4 => SYNTHESIZED_WIRE_313,
		 In_5 => SYNTHESIZED_WIRE_314,
		 In_6 => SYNTHESIZED_WIRE_315,
		 In_7 => SYNTHESIZED_WIRE_316,
		 In_8 => SYNTHESIZED_WIRE_317,
		 Out_0 => SYNTHESIZED_WIRE_340,
		 Out_1 => SYNTHESIZED_WIRE_341,
		 Out_2 => SYNTHESIZED_WIRE_342,
		 Out_3 => SYNTHESIZED_WIRE_343,
		 Out_4 => SYNTHESIZED_WIRE_344,
		 Out_5 => SYNTHESIZED_WIRE_345,
		 Out_6 => SYNTHESIZED_WIRE_346,
		 Out_7 => SYNTHESIZED_WIRE_347,
		 Out_8 => SYNTHESIZED_WIRE_348);


b2v_inst57 : lszd_level3
PORT MAP(MS0 => SYNTHESIZED_WIRE_554,
		 MS1 => SYNTHESIZED_WIRE_555,
		 MS2 => SYNTHESIZED_WIRE_556,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_567,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_566,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_565,
		 NZ_MS => SYNTHESIZED_WIRE_324,
		 NZ_LS => SYNTHESIZED_WIRE_325,
		 P3 => SYNTHESIZED_WIRE_563,
		 P2 => SYNTHESIZED_WIRE_562,
		 P1 => SYNTHESIZED_WIRE_561,
		 P0 => SYNTHESIZED_WIRE_560,
		 NZ => SYNTHESIZED_WIRE_564);


b2v_inst58 : il_level4_new
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_568,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_569,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_570,
		 LSZD_Pos3 => SYNTHESIZED_WIRE_571,
		 LSZD_Pos4 => SYNTHESIZED_WIRE_572,
		 Cout_0 => SYNTHESIZED_WIRE_331,
		 In_0 => SYNTHESIZED_WIRE_573,
		 In_1 => SYNTHESIZED_WIRE_574,
		 In_2 => SYNTHESIZED_WIRE_575,
		 In_3 => SYNTHESIZED_WIRE_576,
		 In_4 => SYNTHESIZED_WIRE_336,
		 In_5 => SYNTHESIZED_WIRE_337,
		 In_6 => SYNTHESIZED_WIRE_338,
		 In_7 => SYNTHESIZED_WIRE_339,
		 In_8 => SYNTHESIZED_WIRE_340,
		 In_9 => SYNTHESIZED_WIRE_341,
		 In_10 => SYNTHESIZED_WIRE_342,
		 In_11 => SYNTHESIZED_WIRE_343,
		 In_12 => SYNTHESIZED_WIRE_344,
		 In_13 => SYNTHESIZED_WIRE_345,
		 In_14 => SYNTHESIZED_WIRE_346,
		 In_15 => SYNTHESIZED_WIRE_347,
		 In_16 => SYNTHESIZED_WIRE_348,
		 Out_0 => SYNTHESIZED_WIRE_24,
		 Out_1 => SYNTHESIZED_WIRE_25,
		 Out_2 => SYNTHESIZED_WIRE_26,
		 Out_3 => SYNTHESIZED_WIRE_27,
		 Out_4 => SYNTHESIZED_WIRE_28,
		 Out_5 => SYNTHESIZED_WIRE_29,
		 Out_6 => SYNTHESIZED_WIRE_30,
		 Out_7 => SYNTHESIZED_WIRE_31,
		 Out_8 => SYNTHESIZED_WIRE_32,
		 Out_9 => SYNTHESIZED_WIRE_33,
		 Out_10 => SYNTHESIZED_WIRE_34,
		 Out_11 => SYNTHESIZED_WIRE_35,
		 Out_12 => SYNTHESIZED_WIRE_36,
		 Out_13 => SYNTHESIZED_WIRE_37,
		 Out_14 => SYNTHESIZED_WIRE_38,
		 Out_15 => SYNTHESIZED_WIRE_39,
		 Out_16 => SYNTHESIZED_WIRE_40);


b2v_inst59 : lszd_level4
PORT MAP(MS0 => SYNTHESIZED_WIRE_560,
		 MS1 => SYNTHESIZED_WIRE_561,
		 MS2 => SYNTHESIZED_WIRE_562,
		 MS3 => SYNTHESIZED_WIRE_563,
		 NZ_MS => SYNTHESIZED_WIRE_564,
		 NZ_LS => SYNTHESIZED_WIRE_536,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_573,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_574,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_575,
		 MSH_LSsumbit_3 => SYNTHESIZED_WIRE_576,
		 P4 => SYNTHESIZED_WIRE_572,
		 P3 => SYNTHESIZED_WIRE_571,
		 P2 => SYNTHESIZED_WIRE_570,
		 P1 => SYNTHESIZED_WIRE_569,
		 P0 => SYNTHESIZED_WIRE_568,
		 NZ => SYNTHESIZED_WIRE_373);


b2v_inst6 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_359,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_360,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_361,
		 Cout_0 => SYNTHESIZED_WIRE_362,
		 In_0 => SYNTHESIZED_WIRE_577,
		 In_1 => SYNTHESIZED_WIRE_578,
		 In_2 => SYNTHESIZED_WIRE_365,
		 In_3 => SYNTHESIZED_WIRE_366,
		 In_4 => SYNTHESIZED_WIRE_367,
		 Out_0 => sum_ALTERA_SYNTHESIZED(4),
		 Out_1 => sum_ALTERA_SYNTHESIZED(5),
		 Out_2 => sum_ALTERA_SYNTHESIZED(6),
		 Out_3 => sum_ALTERA_SYNTHESIZED(7),
		 Out_4 => SYNTHESIZED_WIRE_163);


b2v_inst63 : lszd_level5
PORT MAP(MS0 => SYNTHESIZED_WIRE_568,
		 MS1 => SYNTHESIZED_WIRE_569,
		 MS2 => SYNTHESIZED_WIRE_570,
		 MS3 => SYNTHESIZED_WIRE_571,
		 MS4 => SYNTHESIZED_WIRE_572,
		 NZ_MS => SYNTHESIZED_WIRE_373,
		 NZ_LS => SYNTHESIZED_WIRE_374,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_490,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_491,
		 MSH_LSsumbit_2 => SYNTHESIZED_WIRE_492,
		 MSH_LSsumbit_3 => SYNTHESIZED_WIRE_493,
		 P5 => SYNTHESIZED_WIRE_5,
		 P4 => SYNTHESIZED_WIRE_4,
		 P3 => SYNTHESIZED_WIRE_3,
		 P2 => SYNTHESIZED_WIRE_2,
		 P1 => SYNTHESIZED_WIRE_1,
		 P0 => SYNTHESIZED_WIRE_0,
		 NZ => SYNTHESIZED_WIRE_6);


b2v_inst66 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_579,
		 MS1 => SYNTHESIZED_WIRE_580,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_578,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_577,
		 NZ_MS => SYNTHESIZED_WIRE_383,
		 NZ_LS => SYNTHESIZED_WIRE_384,
		 P2 => SYNTHESIZED_WIRE_361,
		 P1 => SYNTHESIZED_WIRE_360,
		 P0 => SYNTHESIZED_WIRE_359,
		 NZ => SYNTHESIZED_WIRE_279);


b2v_inst67 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_581,
		 MS1 => SYNTHESIZED_WIRE_582,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_583,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_584,
		 NZ_MS => SYNTHESIZED_WIRE_389,
		 NZ_LS => SYNTHESIZED_WIRE_390,
		 P2 => SYNTHESIZED_WIRE_552,
		 P1 => SYNTHESIZED_WIRE_551,
		 P0 => SYNTHESIZED_WIRE_550,
		 NZ => SYNTHESIZED_WIRE_278);


b2v_inst68 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_498,
		 MS1 => SYNTHESIZED_WIRE_499,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_495,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_494,
		 NZ_MS => SYNTHESIZED_WIRE_395,
		 NZ_LS => SYNTHESIZED_WIRE_396,
		 P2 => SYNTHESIZED_WIRE_43,
		 P1 => SYNTHESIZED_WIRE_42,
		 P0 => SYNTHESIZED_WIRE_41,
		 NZ => SYNTHESIZED_WIRE_94);


b2v_inst69 : leaf
PORT MAP(A_1 => a(3),
		 B_1 => b(3),
		 A_0 => a(2),
		 B_0 => b(2),
		 Sum_1p => SYNTHESIZED_WIRE_446,
		 Cout_1p => SYNTHESIZED_WIRE_447,
		 NZ => SYNTHESIZED_WIRE_52,
		 Sum_0 => SYNTHESIZED_WIRE_496,
		 Pos => SYNTHESIZED_WIRE_50);


b2v_inst7 : il_level2
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_550,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_551,
		 LSZD_Pos2 => SYNTHESIZED_WIRE_552,
		 Cout_0 => SYNTHESIZED_WIRE_400,
		 In_0 => SYNTHESIZED_WIRE_584,
		 In_1 => SYNTHESIZED_WIRE_583,
		 In_2 => SYNTHESIZED_WIRE_403,
		 In_3 => SYNTHESIZED_WIRE_404,
		 In_4 => SYNTHESIZED_WIRE_405,
		 Out_0 => SYNTHESIZED_WIRE_168,
		 Out_1 => SYNTHESIZED_WIRE_169,
		 Out_2 => SYNTHESIZED_WIRE_170,
		 Out_3 => SYNTHESIZED_WIRE_171,
		 Out_4 => SYNTHESIZED_WIRE_172);


b2v_inst70 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_585,
		 MS1 => SYNTHESIZED_WIRE_586,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_507,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_506,
		 NZ_MS => SYNTHESIZED_WIRE_410,
		 NZ_LS => SYNTHESIZED_WIRE_411,
		 P2 => SYNTHESIZED_WIRE_505,
		 P1 => SYNTHESIZED_WIRE_504,
		 P0 => SYNTHESIZED_WIRE_503,
		 NZ => SYNTHESIZED_WIRE_93);


b2v_inst71 : leaf
PORT MAP(A_1 => a(19),
		 B_1 => a(19),
		 A_0 => a(18),
		 B_0 => b(18),
		 Sum_1p => SYNTHESIZED_WIRE_452,
		 Cout_1p => SYNTHESIZED_WIRE_453,
		 NZ => SYNTHESIZED_WIRE_66,
		 Sum_0 => SYNTHESIZED_WIRE_501,
		 Pos => SYNTHESIZED_WIRE_64);


b2v_inst72 : leaf
PORT MAP(A_1 => a(17),
		 B_1 => b(17),
		 A_0 => a(16),
		 B_0 => b(16),
		 Sum_1p => SYNTHESIZED_WIRE_524,
		 Cout_1p => SYNTHESIZED_WIRE_450,
		 NZ => SYNTHESIZED_WIRE_67,
		 Sum_0 => SYNTHESIZED_WIRE_523);


b2v_inst73 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_513,
		 MS1 => SYNTHESIZED_WIRE_514,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_512,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_511,
		 NZ_MS => SYNTHESIZED_WIRE_416,
		 NZ_LS => SYNTHESIZED_WIRE_417,
		 P2 => SYNTHESIZED_WIRE_97,
		 P1 => SYNTHESIZED_WIRE_96,
		 P0 => SYNTHESIZED_WIRE_95,
		 NZ => SYNTHESIZED_WIRE_248);


b2v_inst74 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_587,
		 MS1 => SYNTHESIZED_WIRE_588,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_522,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_521,
		 NZ_MS => SYNTHESIZED_WIRE_422,
		 NZ_LS => SYNTHESIZED_WIRE_423,
		 P2 => SYNTHESIZED_WIRE_520,
		 P1 => SYNTHESIZED_WIRE_519,
		 P0 => SYNTHESIZED_WIRE_518,
		 NZ => SYNTHESIZED_WIRE_247);


b2v_inst75 : leaf
PORT MAP(A_1 => a(35),
		 B_1 => b(35),
		 A_0 => a(34),
		 B_0 => b(34),
		 Sum_1p => SYNTHESIZED_WIRE_464,
		 Cout_1p => SYNTHESIZED_WIRE_465,
		 NZ => SYNTHESIZED_WIRE_112,
		 Sum_0 => SYNTHESIZED_WIRE_516,
		 Pos => SYNTHESIZED_WIRE_110);


b2v_inst76 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_546,
		 MS1 => SYNTHESIZED_WIRE_547,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_545,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_544,
		 NZ_MS => SYNTHESIZED_WIRE_428,
		 NZ_LS => SYNTHESIZED_WIRE_429,
		 P2 => SYNTHESIZED_WIRE_251,
		 P1 => SYNTHESIZED_WIRE_250,
		 P0 => SYNTHESIZED_WIRE_249,
		 NZ => SYNTHESIZED_WIRE_325);


b2v_inst77 : lszd_level2_new
PORT MAP(MS0 => SYNTHESIZED_WIRE_589,
		 MS1 => SYNTHESIZED_WIRE_590,
		 MSH_LSsumbit_1 => SYNTHESIZED_WIRE_558,
		 MSH_LSsumbit_0 => SYNTHESIZED_WIRE_557,
		 NZ_MS => SYNTHESIZED_WIRE_434,
		 NZ_LS => SYNTHESIZED_WIRE_435,
		 P2 => SYNTHESIZED_WIRE_556,
		 P1 => SYNTHESIZED_WIRE_555,
		 P0 => SYNTHESIZED_WIRE_554,
		 NZ => SYNTHESIZED_WIRE_324);


b2v_inst773 : leaf_cin
PORT MAP(A_1 => a(1),
		 B_1 => b(1),
		 A_0 => a(0),
		 B_0 => b(0),
		 Cin_init => cin_init,
		 Sum_1p => sum_ALTERA_SYNTHESIZED(1),
		 Cout_1p => SYNTHESIZED_WIRE_444,
		 NZ => SYNTHESIZED_WIRE_53,
		 Sum_0 => sum_ALTERA_SYNTHESIZED(0));


b2v_inst774 : leaf
PORT MAP(A_1 => a(15),
		 B_1 => b(15),
		 A_0 => a(14),
		 B_0 => b(14),
		 Sum_1p => SYNTHESIZED_WIRE_440,
		 Cout_1p => SYNTHESIZED_WIRE_441,
		 NZ => SYNTHESIZED_WIRE_223,
		 Sum_0 => SYNTHESIZED_WIRE_541,
		 Pos => SYNTHESIZED_WIRE_221);


b2v_inst775 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_581,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_582,
		 Cout_0 => SYNTHESIZED_WIRE_438,
		 In_0 => SYNTHESIZED_WIRE_541,
		 In_1 => SYNTHESIZED_WIRE_440,
		 In_2 => SYNTHESIZED_WIRE_441,
		 Out_0 => SYNTHESIZED_WIRE_403,
		 Out_1 => SYNTHESIZED_WIRE_404,
		 Out_2 => SYNTHESIZED_WIRE_405);


b2v_inst776 : leaf
PORT MAP(A_1 => a(5),
		 B_1 => b(5),
		 A_0 => a(4),
		 B_0 => b(4),
		 Sum_1p => SYNTHESIZED_WIRE_578,
		 Cout_1p => SYNTHESIZED_WIRE_486,
		 NZ => SYNTHESIZED_WIRE_220,
		 Sum_0 => SYNTHESIZED_WIRE_577);


b2v_inst777 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_442,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_443,
		 Cout_0 => SYNTHESIZED_WIRE_444,
		 In_0 => SYNTHESIZED_WIRE_496,
		 In_1 => SYNTHESIZED_WIRE_446,
		 In_2 => SYNTHESIZED_WIRE_447,
		 Out_0 => sum_ALTERA_SYNTHESIZED(2),
		 Out_1 => sum_ALTERA_SYNTHESIZED(3),
		 Out_2 => SYNTHESIZED_WIRE_362);


b2v_inst778 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_448,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_449,
		 Cout_0 => SYNTHESIZED_WIRE_450,
		 In_0 => SYNTHESIZED_WIRE_501,
		 In_1 => SYNTHESIZED_WIRE_452,
		 In_2 => SYNTHESIZED_WIRE_453,
		 Out_0 => SYNTHESIZED_WIRE_525,
		 Out_1 => SYNTHESIZED_WIRE_526,
		 Out_2 => SYNTHESIZED_WIRE_44);


b2v_inst779 : leaf
PORT MAP(A_1 => a(21),
		 B_1 => b(21),
		 A_0 => a(20),
		 B_0 => b(20),
		 Sum_1p => SYNTHESIZED_WIRE_495,
		 Cout_1p => SYNTHESIZED_WIRE_60,
		 NZ => SYNTHESIZED_WIRE_228,
		 Sum_0 => SYNTHESIZED_WIRE_494);


b2v_inst78 : leaf
PORT MAP(A_1 => a(51),
		 B_1 => b(51),
		 A_0 => a(50),
		 B_0 => b(50),
		 Sum_1p => SYNTHESIZED_WIRE_476,
		 Cout_1p => SYNTHESIZED_WIRE_477,
		 NZ => SYNTHESIZED_WIRE_266,
		 Sum_0 => SYNTHESIZED_WIRE_549,
		 Pos => SYNTHESIZED_WIRE_264);


b2v_inst780 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_585,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_586,
		 Cout_0 => SYNTHESIZED_WIRE_456,
		 In_0 => SYNTHESIZED_WIRE_542,
		 In_1 => SYNTHESIZED_WIRE_458,
		 In_2 => SYNTHESIZED_WIRE_459,
		 Out_0 => SYNTHESIZED_WIRE_80,
		 Out_1 => SYNTHESIZED_WIRE_81,
		 Out_2 => SYNTHESIZED_WIRE_82);


b2v_inst781 : leaf
PORT MAP(A_1 => a(31),
		 B_1 => b(31),
		 A_0 => a(30),
		 B_0 => b(30),
		 Sum_1p => SYNTHESIZED_WIRE_458,
		 Cout_1p => SYNTHESIZED_WIRE_459,
		 NZ => SYNTHESIZED_WIRE_231,
		 Sum_0 => SYNTHESIZED_WIRE_542,
		 Pos => SYNTHESIZED_WIRE_229);


b2v_inst782 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_460,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_461,
		 Cout_0 => SYNTHESIZED_WIRE_462,
		 In_0 => SYNTHESIZED_WIRE_516,
		 In_1 => SYNTHESIZED_WIRE_464,
		 In_2 => SYNTHESIZED_WIRE_465,
		 Out_0 => SYNTHESIZED_WIRE_492,
		 Out_1 => SYNTHESIZED_WIRE_493,
		 Out_2 => SYNTHESIZED_WIRE_98);


b2v_inst783 : leaf
PORT MAP(A_1 => a(37),
		 B_1 => b(37),
		 A_0 => a(36),
		 B_0 => b(36),
		 Sum_1p => SYNTHESIZED_WIRE_512,
		 Cout_1p => SYNTHESIZED_WIRE_106,
		 NZ => SYNTHESIZED_WIRE_236,
		 Sum_0 => SYNTHESIZED_WIRE_511);


b2v_inst784 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_587,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_588,
		 Cout_0 => SYNTHESIZED_WIRE_468,
		 In_0 => SYNTHESIZED_WIRE_543,
		 In_1 => SYNTHESIZED_WIRE_470,
		 In_2 => SYNTHESIZED_WIRE_471,
		 Out_0 => SYNTHESIZED_WIRE_126,
		 Out_1 => SYNTHESIZED_WIRE_127,
		 Out_2 => SYNTHESIZED_WIRE_128);


b2v_inst785 : leaf
PORT MAP(A_1 => a(47),
		 B_1 => b(47),
		 A_0 => a(46),
		 B_0 => b(46),
		 Sum_1p => SYNTHESIZED_WIRE_470,
		 Cout_1p => SYNTHESIZED_WIRE_471,
		 NZ => SYNTHESIZED_WIRE_239,
		 Sum_0 => SYNTHESIZED_WIRE_543,
		 Pos => SYNTHESIZED_WIRE_237);


b2v_inst787 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_472,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_473,
		 Cout_0 => SYNTHESIZED_WIRE_474,
		 In_0 => SYNTHESIZED_WIRE_549,
		 In_1 => SYNTHESIZED_WIRE_476,
		 In_2 => SYNTHESIZED_WIRE_477,
		 Out_0 => SYNTHESIZED_WIRE_575,
		 Out_1 => SYNTHESIZED_WIRE_576,
		 Out_2 => SYNTHESIZED_WIRE_252);


b2v_inst788 : leaf
PORT MAP(A_1 => a(53),
		 B_1 => b(53),
		 A_0 => a(52),
		 B_0 => b(52),
		 Sum_1p => SYNTHESIZED_WIRE_545,
		 Cout_1p => SYNTHESIZED_WIRE_260,
		 NZ => SYNTHESIZED_WIRE_271,
		 Sum_0 => SYNTHESIZED_WIRE_544);


b2v_inst789 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_589,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_590,
		 Cout_0 => SYNTHESIZED_WIRE_480,
		 In_0 => SYNTHESIZED_WIRE_559,
		 In_1 => SYNTHESIZED_WIRE_482,
		 In_2 => SYNTHESIZED_WIRE_483,
		 Out_0 => SYNTHESIZED_WIRE_292,
		 Out_1 => SYNTHESIZED_WIRE_293,
		 Out_2 => SYNTHESIZED_WIRE_294);


b2v_inst79 : leaf
PORT MAP(A_1 => a(49),
		 B_1 => b(49),
		 A_0 => a(48),
		 B_0 => b(48),
		 Sum_1p => SYNTHESIZED_WIRE_574,
		 Cout_1p => SYNTHESIZED_WIRE_474,
		 NZ => SYNTHESIZED_WIRE_267,
		 Sum_0 => SYNTHESIZED_WIRE_573);


b2v_inst790 : leaf
PORT MAP(A_1 => a(63),
		 B_1 => b(63),
		 A_0 => a(62),
		 B_0 => b(62),
		 Sum_1p => SYNTHESIZED_WIRE_482,
		 Cout_1p => SYNTHESIZED_WIRE_483,
		 NZ => SYNTHESIZED_WIRE_301,
		 Sum_0 => SYNTHESIZED_WIRE_559,
		 Pos => SYNTHESIZED_WIRE_299);


b2v_inst8 : il_level1s
PORT MAP(LSZD_Pos0 => SYNTHESIZED_WIRE_579,
		 LSZD_Pos1 => SYNTHESIZED_WIRE_580,
		 Cout_0 => SYNTHESIZED_WIRE_486,
		 In_0 => SYNTHESIZED_WIRE_540,
		 In_1 => SYNTHESIZED_WIRE_488,
		 In_2 => SYNTHESIZED_WIRE_489,
		 Out_0 => SYNTHESIZED_WIRE_365,
		 Out_1 => SYNTHESIZED_WIRE_366,
		 Out_2 => SYNTHESIZED_WIRE_367);


b2v_inst80 : leaf
PORT MAP(A_1 => a(33),
		 B_1 => b(33),
		 A_0 => a(32),
		 B_0 => b(32),
		 Sum_1p => SYNTHESIZED_WIRE_491,
		 Cout_1p => SYNTHESIZED_WIRE_462,
		 NZ => SYNTHESIZED_WIRE_113,
		 Sum_0 => SYNTHESIZED_WIRE_490);


b2v_inst9 : leaf
PORT MAP(A_1 => a(7),
		 B_1 => b(7),
		 A_0 => a(6),
		 B_0 => b(6),
		 Sum_1p => SYNTHESIZED_WIRE_488,
		 Cout_1p => SYNTHESIZED_WIRE_489,
		 NZ => SYNTHESIZED_WIRE_219,
		 Sum_0 => SYNTHESIZED_WIRE_540,
		 Pos => SYNTHESIZED_WIRE_217);

sum <= sum_ALTERA_SYNTHESIZED;

END bdf_type;